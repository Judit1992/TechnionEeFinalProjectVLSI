/**
 *-----------------------------------------------------
 * Module Name: 	ga_init_pop
 * Author 	  :		Judit Ben Ami , May Buzaglo
 * Date		  : 	September 23, 2021
 *-----------------------------------------------------
 *
 * Module Description:
 * =================================
 *
 *
 */
 

module ga_crossover_find_thresholds #(
	`include "ga_params.const"
	) ( 
	//***********************************
	// Cnfg
	//***********************************
	//inputs
	input [FIT_SCORE_W-1:0]			cnfg_max_fit_socre,	
	//***********************************
	// Data IF: GA_CROSSOVER <-> SELF
	//***********************************
	//outputs
	output logic [FIT_SCORE_W-1:0]		thresh_ary [0:DATA_W-1] //1 thresh per bit
	);


// =========================================================================
// local parameters and ints
// =========================================================================
genvar gv0;


// =========================================================================
// signals decleration
// =========================================================================


// #########################################################################
// #########################################################################
// ------------------------- MODULE LOGIC ----------------------------------
// #########################################################################
// #########################################################################

assign thresh_ary[0] = { {(FIT_SCORE_INT_W-1){1'b0}} , 1'b1 , {FIT_SCORE_FRACT_W{1'b0}} } >> (DATA_W-1); //2^-(DATA_W-1)
generate 
	for (gv0=1;gv0<DATA_W;gv0++)
		begin: CREATE_THRESH_LOOP
		assign thresh_ary[gv0] = cnfg_max_fit_socre >> (DATA_W-gv0);
		end
endgenerate


endmodule



